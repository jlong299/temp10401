
module ROM_sin_dct_vecRot (
	address,
	clock,
	q);	

	input	[10:0]	address;
	input		clock;
	output	[17:0]	q;
endmodule
